��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  !	G    Alarma      �  )^7    Bomba de Entrada      �  �p�    Bomba de Salida      �  �� ��     Sensor C      �  q� ��     Sensor B      �  � G�     Sensor A                    ��� 	 CLogicOut�� 	 CTerminal   H5I              @            4@DP          ��    ��  8(M)               �            L \0           ��    �� 	 CRailThru�  �`�u       d       @          �  �d�y     
         @            �b�v        ����    ��  � �5       d       @          �  �$�9              @            �"�6        ����    ��  CAND�  � �!               �          �  �0�1              @          �  �(�)               �            ��4           ��    ��  @ U                          �  @U                          �  l�	               �            T�l     "      ��    ��  @�U�     	 	       @            T�d�     &     ��    ��  CNAND�   ��               �          �   ��              @          �  ,�A�     	         @            �,�     )      ��    '��  ����              @          �  ����              @          �  ����               �            ����     -      ��    '��  0�E�              @          �  0�E�                          �  \�q�              @            D�\�     1      ��    '��  0�E�                          �  0�E�                          �  \�q�              @            D�\�     5      ��    ��  CNOR�  8@MA                          �  8PMQ                          �  dHyI              @            L<dT     :      ��    ��  ��-       d       @          �  ��1              @            ��.    >    ����    ��  �0�E       d                   �  �4�I                            �2�F    A    ����    ��  ��-       d                   �  ��1                            ��.    D    ����    ��  @0AE       d                   �  @4AI                            <2DF    G    ����    ��  @0AE       d                   �  @4AI                            <2DF    J    ����    ��  @A-       d                   �  @A1                            <D.    M    ����    ��  CLogicIn�� 	 CLatchKey  �� �     P   �  ��              @            �� �    S   ����     ��  ��              @            �� �    U     ��    O�Q�  x� �      V   �  ��                            �� �    X    ����     ��  pq                            h� x    Z      ��    O�Q�  (� 8      [   �  @A                            <� D    ]    ����     ��   !                            � (    _      ��                  ���  CWire  xH!I      a�  �(9)      a�  �H�a       a�  �8�I       a�  �HI      a�   0I       a�   0�1      a��� 
 CCrossOver  ��      j�  ���      j�  ����        ���!       a�j�  ��        �A      a�j�  ���      j�  ���        @ A      a�j�  ����        ��1�      a�  ��1�      a�j�  ����      j�  ����        @�1�      a�  � �!      a�  ��!       a�  ��1       a�j�  ���        ���       a�  @ A1       a�  @�A       a�  @`A�       a�j�  �<�D      j�  �L�T      j�  ����        �0��       a�  p�q�       a�  p��      a�   ��       a�  ���      a�j�  ����        �P��       a�  ����       a�  ����      a�  ����       a�  p���      a�  0�1�       a�j�  �<�D        �0�Q       a�j�  �L�T        �P9Q      a�  @HAa       a�  @`Qa      a�  P@Qa       a�j�  �<�D      j�  �<�D        P@9A      a�  ��      a�   A      a�  p�                    �                             b   c  d      i    e  y   h      c " p " # n # $ $ z & + & ) � ) * � * + + & - � - . � . / / � 1 u 1 2 s 2 3 3 � 5 � 5 6 � 6 7 7 � : � : ; � ; < < b S > ? ? � { A B B   X D E E � ~ G H H   N J K K � ] M N N J S S � U U � X X � Z Z � ] ] � _ _ � <     e   f d g h f g  i o i q i t �  n k { # p l p } ~ " s m | 2 i 1 v � v �  5 z  $ y | A | r � n  G � p � v � � � � � x ? � � 3 � * � ) / � � w � s � u � . � - 7 � v 6 � � E � � � � ; K � � � � � � � � � � : U > _ M Z D             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 